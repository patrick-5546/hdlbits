module top_module (
    input  in,
    output out
);

  // bitwise-NOT: ~
  // logical-NOT: !
  assign out = ~in;

endmodule
